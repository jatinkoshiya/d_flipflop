module d_fp 
  begin

  end
endmodule
